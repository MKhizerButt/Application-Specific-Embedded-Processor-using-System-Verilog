// alucodes or ALUfunc[1:0]
`define RA    2'b00
`define RMUL  2'b01
`define RADD  2'b10
`define RSUB  2'b11  